/*+++++++++++++++++++++++++++++++++++
author:qqyk
++ 
++ 
+++++++++++++++++++++++++++++++++++++*/
module gf_mul_8 (
	input wire [7:0] a,
	input wire [7:0] b,
	output wire [7:0] out
	);


	assign out[0] = (a[0]^b[0])^(a[1]^b[7])^(a[2]^b[6])^(a[3]^b[5])^(a[4]^b[4])^(a[5]^b[3])^(a[5]^b[7])^(a[6]^b[2])^(a[6]^b[6])^(a[6]^b[7])^(a[7]^b[1])^(a[7]^b[5])^(a[7]^b[6])^(a[7]^b[7]);
	assign out[1] = (a[0]^b[1])^(a[1]^b[0])^(a[2]^b[7])^(a[3]^b[6])^(a[4]^b[5])^(a[5]^b[4])^(a[6]^b[3])^(a[6]^b[7])^(a[7]^b[2])^(a[7]^b[6])^(a[7]^b[7]);
	assign out[2] = (a[0]^b[2])^(a[1]^b[1])^(a[1]^b[7])^(a[2]^b[0])^(a[2]^b[6])^(a[3]^b[5])^(a[3]^b[7])^(a[4]^b[4])^(a[4]^b[6])^(a[5]^b[3])^(a[5]^b[5])^(a[5]^b[7])^(a[6]^b[2])^(a[6]^b[4])^(a[6]^b[6])^(a[6]^b[7])^(a[7]^b[1])^(a[7]^b[3])^(a[7]^b[5])^(a[7]^b[6]);
	assign out[3] = (a[0]^b[3])^(a[1]^b[2])^(a[1]^b[7])^(a[2]^b[1])^(a[2]^b[6])^(a[2]^b[7])^(a[3]^b[0])^(a[3]^b[5])^(a[3]^b[6])^(a[4]^b[4])^(a[4]^b[5])^(a[4]^b[7])^(a[5]^b[3])^(a[5]^b[4])^(a[5]^b[6])^(a[5]^b[7])^(a[6]^b[2])^(a[6]^b[3])^(a[6]^b[5])^(a[6]^b[6])^(a[7]^b[1])^(a[7]^b[2])^(a[7]^b[4])^(a[7]^b[5]);
	assign out[4] = (a[0]^b[4])^(a[1]^b[3])^(a[1]^b[7])^(a[2]^b[2])^(a[2]^b[6])^(a[2]^b[7])^(a[3]^b[1])^(a[3]^b[5])^(a[3]^b[6])^(a[3]^b[7])^(a[4]^b[0])^(a[4]^b[4])^(a[4]^b[5])^(a[4]^b[6])^(a[5]^b[3])^(a[5]^b[4])^(a[5]^b[5])^(a[6]^b[2])^(a[6]^b[3])^(a[6]^b[4])^(a[7]^b[1])^(a[7]^b[2])^(a[7]^b[3])^(a[7]^b[7]);
	assign out[5] = (a[0]^b[5])^(a[1]^b[4])^(a[2]^b[3])^(a[2]^b[7])^(a[3]^b[2])^(a[3]^b[6])^(a[3]^b[7])^(a[4]^b[1])^(a[4]^b[5])^(a[4]^b[6])^(a[4]^b[7])^(a[5]^b[0])^(a[5]^b[4])^(a[5]^b[5])^(a[5]^b[6])^(a[6]^b[3])^(a[6]^b[4])^(a[6]^b[5])^(a[7]^b[2])^(a[7]^b[3])^(a[7]^b[4]);
	assign out[6] = (a[0]^b[6])^(a[1]^b[5])^(a[2]^b[4])^(a[3]^b[3])^(a[3]^b[7])^(a[4]^b[2])^(a[4]^b[6])^(a[4]^b[7])^(a[5]^b[1])^(a[5]^b[5])^(a[5]^b[6])^(a[5]^b[7])^(a[6]^b[0])^(a[6]^b[4])^(a[6]^b[5])^(a[6]^b[6])^(a[7]^b[3])^(a[7]^b[4])^(a[7]^b[5]);
	assign out[7] = (a[0]^b[7])^(a[1]^b[6])^(a[2]^b[5])^(a[3]^b[4])^(a[4]^b[3])^(a[4]^b[7])^(a[5]^b[2])^(a[5]^b[6])^(a[5]^b[7])^(a[6]^b[1])^(a[6]^b[5])^(a[6]^b[6])^(a[6]^b[7])^(a[7]^b[0])^(a[7]^b[4])^(a[7]^b[5])^(a[7]^b[6]);
endmodule
